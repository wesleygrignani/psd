library ieee;
use ieee.std_logic_1164.all;

package filter_pkg is

  constant KERNEL_SIZE : integer := 3;
  constant IMG_WIDTH   : integer := 256;

end package filter_pkg;