library ieee;
use ieee.std_logic_1164.all;

entity encoder is
  port (
  );
end entity;